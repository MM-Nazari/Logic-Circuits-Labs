`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:31:12 11/30/2021 
// Design Name: 
// Module Name:    Lab8 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module alu(y , A , B ,s );
input [1:0] A , B ;
input [3:0] y ; 
input [1:0] s ;
wire [3:0] w3 ;
wire [2:0] w2 ;
wire [1:0] w1,w0 ;
assign w3 = A*B;
assign w2 = A + B;
assign w1 = ~(A&B);
assign w0 = ~A;

assign y = s[1] ? (s[0] ? w3 : {1'b0,w2} ) : ( s[0] ? {2'b00,w1} : {2'b00,w0});

endmodule
module tb_alu ();


reg [1:0] A;
reg [1:0] B;
reg [1:0] sel;
wire [3:0] Y;

	alu test_alu (Y,A,B,sel);

	initial 
		begin
		A <= 2'b00;
		B <= 2'b00;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b00;
		B <= 2'b01;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b01;
		B <= 2'b00;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b01;
		B <= 2'b01;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b00;
		B <= 2'b10;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b00;
		B <= 2'b11;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b01;
		B <= 2'b10;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b01;
		B <= 2'b11;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b10;
		B <= 2'b00;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b10;
		B <= 2'b01;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b11;
		B <= 2'b00;
		sel <= 2'b00;
		# 10;

		A <= 2'b11;
		B <= 2'b01;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b10;
		B <= 2'b10;
		sel <= 2'b00;
		# 10;

		A <= 2'b10;
		B <= 2'b11;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b11;
		B <= 2'b10;
		sel <= 2'b00;
		# 10;
			
		A <= 2'b11;
		B <= 2'b11;
		sel <= 2'b00;
		# 10;
		
		//******************************************************
		
		A <= 2'b00;
		B <= 2'b00;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b00;
		B <= 2'b01;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b01;
		B <= 2'b00;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b01;
		B <= 2'b01;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b00;
		B <= 2'b10;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b00;
		B <= 2'b11;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b01;
		B <= 2'b10;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b01;
		B <= 2'b11;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b10;
		B <= 2'b00;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b10;
		B <= 2'b01;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b11;
		B <= 2'b00;
		sel <= 2'b01;
		# 10;

		A <= 2'b11;
		B <= 2'b01;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b10;
		B <= 2'b10;
		sel <= 2'b01;
		# 10;

		A <= 2'b10;
		B <= 2'b11;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b11;
		B <= 2'b10;
		sel <= 2'b01;
		# 10;
			
		A <= 2'b11;
		B <= 2'b11;
		sel <= 2'b01;
		# 10;
		//*********************************
		
		A <= 2'b00;
		B <= 2'b00;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b00;
		B <= 2'b01;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b01;
		B <= 2'b00;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b01;
		B <= 2'b01;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b00;
		B <= 2'b10;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b00;
		B <= 2'b11;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b01;
		B <= 2'b10;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b01;
		B <= 2'b11;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b10;
		B <= 2'b00;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b10;
		B <= 2'b01;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b11;
		B <= 2'b00;
		sel <= 2'b10;
		# 10;

		A <= 2'b11;
		B <= 2'b01;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b10;
		B <= 2'b10;
		sel <= 2'b10;
		# 10;

		A <= 2'b10;
		B <= 2'b11;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b11;
		B <= 2'b10;
		sel <= 2'b10;
		# 10;
			
		A <= 2'b11;
		B <= 2'b11;
		sel <= 2'b10;
		# 10;
		
		//***********************************************
		A <= 2'b00;
		B <= 2'b00;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b00;
		B <= 2'b01;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b01;
		B <= 2'b00;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b01;
		B <= 2'b01;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b00;
		B <= 2'b10;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b00;
		B <= 2'b11;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b01;
		B <= 2'b10;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b01;
		B <= 2'b11;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b10;
		B <= 2'b00;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b10;
		B <= 2'b01;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b11;
		B <= 2'b00;
		sel <= 2'b11;
		# 10;

		A <= 2'b11;
		B <= 2'b01;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b10;
		B <= 2'b10;
		sel <= 2'b11;
		# 10;

		A <= 2'b10;
		B <= 2'b11;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b11;
		B <= 2'b10;
		sel <= 2'b11;
		# 10;
			
		A <= 2'b11;
		B <= 2'b11;
		sel <= 2'b11;
		# 10;
		
	
	end

endmodule

